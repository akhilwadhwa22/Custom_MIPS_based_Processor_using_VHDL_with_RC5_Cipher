library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

PACKAGE state_pkg IS
    TYPE s_type is (PKG,KG,IRC,IRD,ENCRYPT,DECRYPT);
END state_pkg;